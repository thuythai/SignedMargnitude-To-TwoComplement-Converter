//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "moodle.v"
//: property showSwitchNets = 0
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w7;    //: /sn:0 {0}(-141,-123)(-131,-123)(-131,23)(-28,23){1}
reg w0;    //: /sn:0 {0}(-28,-7)(-30,-7)(-30,-31)(40,-31)(40,-123)(25,-123){1}
reg w2;    //: /sn:0 {0}(-28,2)(-39,2)(-39,-52)(-29,-52)(-29,-123)(-33,-123){1}
reg w5;    //: /sn:0 {0}(-85,-123)(-75,-123)(-75,13)(-28,13){1}
wire w6;    //: /sn:0 {0}(51,29)(70,29)(70,52)(145,52){1}
//: {2}(149,52)(305,52)(305,175)(346,175){3}
//: {4}(147,50)(147,-37){5}
wire w51;    //: /sn:0 {0}(51,-7)(91,-7)(91,21)(273,21){1}
//: {2}(277,21)(321,21)(321,145)(346,145){3}
//: {4}(275,19)(275,-38){5}
wire w34;    //: /sn:0 {0}(51,2)(88,2)(88,30)(248,30){1}
//: {2}(252,30)(316,30)(316,154)(346,154){3}
//: {4}(250,28)(250,-38){5}
wire w20;    //: /sn:0 {0}(513,115)(513,165)(425,165){1}
wire w17;    //: /sn:0 {0}(598,112)(598,145)(425,145){1}
wire w11;    //: /sn:0 {0}(464,118)(464,181)(425,181){1}
wire w13;    //: /sn:0 {0}(558,114)(558,154)(425,154){1}
wire w9;    //: /sn:0 {0}(51,13)(81,13)(81,41)(191,41){1}
//: {2}(195,41)(311,41)(311,165)(346,165){3}
//: {4}(193,39)(193,-37){5}
//: enddecls

  //: LED g8 (w9) @(193,-44) /sn:0 /w:[ 5 ] /type:0
  //: SWITCH g4 (w2) @(-50,-123) /sn:0 /w:[ 1 ] /st:1 /dn:0
  twosComp g3 (.I0(w0), .I1(w2), .I2(w5), .I3(w7), .O0(w51), .O1(w34), .O2(w9), .O3(w6));   //: @(-27, -17) /sz:(77, 96) /sn:0 /p:[ Li0>0 Li1>0 Li2>1 Li3>1 Ro0<0 Ro1<0 Ro2<0 Ro3<0 ]
  //: comment g1 @(370,-166) /sn:0
  //: /line:"Signed    |  Signed Two's"
  //: /line:"Magnitude |   Complement"
  //: /line:"0111      |   0111"
  //: /line:"0110      |   0110"
  //: /line:"0101      |   0101"
  //: /line:"0100      |   0100"
  //: /line:"0011      |   0011"
  //: /line:"0010      |   0010"
  //: /line:"0001      |   0001"
  //: /line:"0000      |   0000"
  //: /line:""
  //: /line:"1000      |   0000"
  //: /line:"1001      |   1111"
  //: /line:"1010      |   1110"
  //: /line:"1011      |   1101"
  //: /line:"1100      |   1100"
  //: /line:"1101      |   1011"
  //: /line:"1110      |   1010"
  //: /line:"1111      |   1001"
  //: /line:"          "
  //: /line:""
  //: /end
  //: LED g16 (w13) @(558,107) /sn:0 /w:[ 0 ] /type:0
  //: joint g11 (w9) @(193, 41) /w:[ 2 4 1 -1 ]
  //: joint g10 (w6) @(147, 52) /w:[ 2 4 1 -1 ]
  //: joint g19 (w51) @(275, 21) /w:[ 2 4 1 -1 ]
  //: SWITCH g6 (w5) @(-102,-123) /sn:0 /w:[ 0 ] /st:1 /dn:0
  //: LED g7 (w6) @(147,-44) /sn:0 /w:[ 5 ] /type:0
  //: LED g9 (w51) @(275,-45) /sn:0 /w:[ 5 ] /type:0
  //: LED g15 (w17) @(598,105) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g20 (w0) @(8,-123) /sn:0 /w:[ 1 ] /st:1 /dn:0
  //: LED g17 (w20) @(513,108) /sn:0 /w:[ 0 ] /type:0
  //: LED g5 (w34) @(250,-45) /sn:0 /w:[ 5 ] /type:0
  //: SWITCH g21 (w7) @(-158,-123) /sn:0 /w:[ 0 ] /st:0 /dn:0
  twosComp g0 (.I0(w51), .I1(w34), .I2(w9), .I3(w6), .O0(w17), .O1(w13), .O2(w20), .O3(w11));   //: @(347, 135) /sz:(77, 96) /sn:0 /p:[ Li0>3 Li1>3 Li2>3 Li3>3 Ro0<1 Ro1<1 Ro2<1 Ro3<1 ]
  //: LED g18 (w11) @(464,111) /sn:0 /w:[ 0 ] /type:0
  //: joint g12 (w34) @(250, 30) /w:[ 2 4 1 -1 ]

endmodule
//: /netlistEnd

//: /netlistBegin newTwoComp
module newTwoComp();
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
//: enddecls


endmodule
//: /netlistEnd

//: /netlistBegin twosComp
module twosComp(O3, I2, I1, O0, O1, I3, O2, I0);
//: interface  /sz:(77, 96) /bd:[ Li0>I0(10/96) Li1>I1(19/96) Li2>I2(30/96) Li3>I3(40/96) Ro0<O0(10/96) Ro1<O1(19/96) Ro2<O2(30/96) Ro3<O3(46/96) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input I2;    //: /sn:0 {0}(385,138)(263,138)(263,157)(44,157){1}
//: {2}(42,155)(42,5){3}
//: {4}(44,3)(377,3){5}
//: {6}(42,1)(42,-36)(376,-36){7}
//: {8}(42,159)(42,218){9}
//: {10}(44,220)(305,220)(305,211)(468,211){11}
//: {12}(42,222)(42,396)(14,396){13}
input I1;    //: /sn:0 {0}(15,441)(145,441)(145,319){1}
//: {2}(147,317)(355,317){3}
//: {4}(143,317)(142,317)(142,246){5}
//: {6}(144,244)(423,244){7}
//: {8}(142,242)(142,232){9}
//: {10}(144,230)(321,230)(321,216)(468,216){11}
//: {12}(142,228)(142,171){13}
//: {14}(144,169)(210,169){15}
//: {16}(142,167)(142,-31)(376,-31){17}
output O3;    //: /sn:0 {0}(581,-79)(681,-79){1}
input I0;    //: /sn:0 {0}(468,221)(339,221)(339,501){1}
//: {2}(341,503)(551,503)(551,494){3}
//: {4}(553,492)(594,492)(594,493)(615,493){5}
//: {6}(551,490)(551,478)(600,478)(600,488)(615,488){7}
//: {8}(337,503)(243,503){9}
//: {10}(241,501)(241,322)(355,322){11}
//: {12}(239,503)(193,503){13}
//: {14}(191,501)(191,174)(210,174){15}
//: {16}(189,503)(166,503){17}
//: {18}(164,501)(164,-26)(376,-26){19}
//: {20}(162,503)(12,503){21}
output O2;    //: /sn:0 {0}(596,6)(716,6){1}
output O1;    //: /sn:0 {0}(712,245)(608,245){1}
output O0;    //: /sn:0 {0}(636,491)(745,491){1}
input I3;    //: /sn:0 {0}(468,206)(20,206){1}
//: {2}(18,204)(18,135){3}
//: {4}(20,133)(385,133){5}
//: {6}(18,131)(18,0){7}
//: {8}(20,-2)(377,-2){9}
//: {10}(18,-4)(18,-82)(560,-82){11}
//: {12}(18,208)(18,237){13}
//: {14}(20,239)(423,239){15}
//: {16}(18,241)(18,287){17}
//: {18}(20,289)(428,289){19}
//: {20}(18,291)(18,367)(12,367){21}
wire w7;    //: /sn:0 {0}(231,172)(287,172)(287,143)(385,143){1}
wire w4;    //: /sn:0 {0}(489,213)(564,213)(564,11)(575,11){1}
wire w0;    //: /sn:0 {0}(398,1)(575,1){1}
wire w1;    //: /sn:0 {0}(397,-31)(550,-31)(550,-77)(560,-77){1}
wire w8;    //: /sn:0 {0}(449,292)(576,292)(576,247)(587,247){1}
wire w2;    //: /sn:0 {0}(575,6)(502,6)(502,138)(406,138){1}
wire w10;    //: /sn:0 {0}(376,320)(421,320)(421,294)(428,294){1}
wire w5;    //: /sn:0 {0}(444,242)(587,242){1}
//: enddecls

  //: OUT g4 (O3) @(678,-79) /sn:0 /w:[ 1 ]
  _GGOR2 #(6) g8 (.I0(w5), .I1(w8), .Z(O1));   //: @(598,245) /sn:0 /w:[ 1 1 1 ]
  //: joint g13 (I2) @(42, 3) /w:[ 4 6 -1 3 ]
  //: joint g34 (I0) @(191, 503) /w:[ 13 14 16 -1 ]
  _GGAND2 #(6) g3 (.I0(I0), .I1(I0), .Z(O0));   //: @(626,491) /sn:0 /w:[ 7 5 0 ]
  //: IN g2 (I2) @(12,396) /sn:0 /w:[ 13 ]
  //: IN g1 (I1) @(12,441) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g11 (.I0(!I3), .I1(I2), .Z(w0));   //: @(388,1) /sn:0 /w:[ 9 5 0 ]
  _GGOR2 #(6) g16 (.I0(I1), .I1(I0), .Z(w7));   //: @(221,172) /sn:0 /w:[ 15 15 0 ]
  _GGOR3 #(8) g10 (.I0(w0), .I1(w2), .I2(w4), .Z(O2));   //: @(586,6) /sn:0 /w:[ 1 0 1 0 ]
  //: joint g28 (I0) @(164, 503) /w:[ 17 18 20 -1 ]
  //: OUT g32 (O0) @(742,491) /sn:0 /w:[ 1 ]
  //: joint g19 (I3) @(18, 206) /w:[ 1 2 -1 12 ]
  _GGAND2 #(6) g27 (.I0(I3), .I1(w10), .Z(w8));   //: @(439,292) /sn:0 /w:[ 19 1 0 ]
  //: OUT g6 (O1) @(709,245) /sn:0 /w:[ 0 ]
  _GGOR3 #(8) g9 (.I0(I2), .I1(I1), .I2(I0), .Z(w1));   //: @(387,-31) /sn:0 /w:[ 7 17 19 0 ]
  //: joint g7 (I0) @(551, 492) /w:[ 4 6 -1 3 ]
  //: IN g31 (I3) @(10,367) /sn:0 /w:[ 21 ]
  //: joint g15 (I2) @(42, 157) /w:[ 1 2 -1 8 ]
  //: joint g20 (I2) @(42, 220) /w:[ 10 9 -1 12 ]
  //: joint g17 (I1) @(142, 169) /w:[ 14 16 -1 13 ]
  //: joint g25 (I3) @(18, 239) /w:[ 14 13 -1 16 ]
  _GGXOR2 #(8) g29 (.I0(I1), .I1(I0), .Z(w10));   //: @(366,320) /sn:0 /w:[ 3 11 0 ]
  //: OUT g5 (O2) @(713,6) /sn:0 /w:[ 1 ]
  _GGAND3 #(8) g14 (.I0(I3), .I1(!I2), .I2(w7), .Z(w2));   //: @(396,138) /sn:0 /w:[ 5 0 1 1 ]
  //: joint g21 (I1) @(142, 230) /w:[ 10 12 -1 9 ]
  //: joint g24 (I3) @(18, 133) /w:[ 4 6 -1 3 ]
  //: joint g36 (I0) @(339, 503) /w:[ 2 1 8 -1 ]
  _GGAND2 #(6) g23 (.I0(!I3), .I1(I1), .Z(w5));   //: @(434,242) /sn:0 /w:[ 15 7 0 ]
  //: IN g0 (I0) @(10,503) /sn:0 /w:[ 21 ]
  _GGAND2 #(6) g22 (.I0(I3), .I1(w1), .Z(O3));   //: @(571,-79) /sn:0 /w:[ 11 1 0 ]
  //: joint g26 (I1) @(142, 244) /w:[ 6 8 -1 5 ]
  //: joint g35 (I0) @(241, 503) /w:[ 9 10 12 -1 ]
  _GGAND4 #(10) g18 (.I0(I3), .I1(I2), .I2(!I1), .I3(!I0), .Z(w4));   //: @(479,213) /sn:0 /w:[ 0 11 11 0 0 ]
  //: joint g12 (I3) @(18, -2) /w:[ 8 10 -1 7 ]
  //: joint g33 (I3) @(18, 289) /w:[ 18 17 -1 20 ]
  //: joint g30 (I1) @(145, 317) /w:[ 2 -1 4 1 ]

endmodule
//: /netlistEnd

